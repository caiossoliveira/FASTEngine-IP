LIBRARY IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.numeric_std.all;

use work.fast_engine_types.all;

ENTITY test_FASTEngine IS
END ENTITY;

ARCHITECTURE test_FASTEngine OF test_FASTEngine IS
  COMPONENT FASTEngine IS
    port (
		clk: in STD_LOGIC;
		reset: in STD_LOGIC;
		enable: in STD_LOGIC;

        FASTByte_in: in STD_LOGIC_VECTOR (7 downto 0);
		read_in: in STD_LOGIC;

		startOfMachine_out: out STD_LOGIC;
		reading_out: out STD_LOGIC;

		type_out : out STD_LOGIC;
        updateAction_out : out STD_LOGIC_VECTOR(6 downto 0);
		position_out : out STD_LOGIC_VECTOR(3 downto 0);
		size_out : out STD_LOGIC_VECTOR(63 downto 0);
		exp_out : out STD_LOGIC_VECTOR(31 downto 0);
		man_out : out STD_LOGIC_VECTOR(63 downto 0);

        ready_out : out STD_LOGIC
	);
  END COMPONENT;

  SIGNAL counter : INTEGER;
  SIGNAL sig_aux_counter : STD_LOGIC;
  
  SIGNAL sig_clk    : STD_LOGIC := '0';
  SIGNAL sig_reset  : STD_LOGIC;
  SIGNAL sig_msg_in : STD_LOGIC_VECTOR (7 DOWNTO 0);
  SIGNAL sig_enable : STD_LOGIC := '0';

  SIGNAL sig_read   : STD_LOGIC;
  SIGNAL sig_startOfMachine :   STD_LOGIC;
  SIGNAL sig_reading    : STD_LOGIC := '0';

  SIGNAL sig_type_out : STD_LOGIC;
  SIGNAL sig_updateAction_out : STD_LOGIC_VECTOR(6 downto 0);
  SIGNAL sig_position_out : STD_LOGIC_VECTOR(3 downto 0);
  SIGNAL sig_size_out : STD_LOGIC_VECTOR(63 downto 0);
  SIGNAL sig_exp_out : STD_LOGIC_VECTOR(31 downto 0);
  SIGNAL sig_man_out : STD_LOGIC_VECTOR(63 downto 0);

  SIGNAL sig_ready_out : STD_LOGIC;

  SIGNAL sig_test_out : STD_LOGIC_VECTOR(7 downto 0);

  -- FASTMem signals declarations
  signal sl_enableFASTMem: STD_LOGIC;
  signal mem_counter: INTEGER := 0;
  signal FASTByte: STD_LOGIC_VECTOR (7 downto 0);

  -- book signals declarations
  signal bidOrderDepthBook_size : POSITION_TYPE_SIZE(0 to 9) := (OTHERS => X"0000000000000000");
  signal bidOrderDepthBook_px_exp : POSITION_TYPE_PX_EXP(0 to 9) := (OTHERS => X"00000000");
  signal bidOrderDepthBook_px_man : POSITION_TYPE_PX_MAN(0 to 9) := (OTHERS => X"FFFFFFFFFFFFFFFF");

  signal offerOrderDepthBook_size : POSITION_TYPE_SIZE(0 to 9) := (OTHERS => X"0000000000000000");
  signal offerOrderDepthBook_px_exp : POSITION_TYPE_PX_EXP(0 to 9) := (OTHERS => X"00000000");
  signal offerOrderDepthBook_px_man : POSITION_TYPE_PX_MAN(0 to 9) := (OTHERS => X"FFFFFFFFFFFFFFFF");

  -- SYMBOLIC ENCODED state machine: FASTMem
  type FASTMem_type is (
      Start, writeByte
  );
 -- attribute ENUM_ENCODING of FASTMem_type: type is ... -- enum_encoding attribute is not supported for symbolic encoding

signal FASTMem, NextState_FASTMem: FASTMem_type;

-- Declarations of pre-registered internal signals
--signal int_msg_out, next_msg_out: STD_LOGIC_VECTOR (7 downto 0);
signal next_mem_counter: INTEGER := 0;
--signal next_mem_out: STD_LOGIC_VECTOR (7 downto 0);
--signal next_FASTByte : STD_LOGIC_VECTOR (7 downto 0);
signal next_sig_msg_in : STD_LOGIC_VECTOR( 7 DOWNTO 0);
--signal next_read: STD_LOGIC;
--signal next_sig_read : STD_LOGIC;
--signal next_reading: STD_LOGIC;
--signal next_startOfMachine: STD_LOGIC;


BEGIN
    fe  : FASTEngine  PORT MAP (clk => sig_clk, reset => sig_reset, FASTByte_in => sig_msg_in, enable => sig_enable,
                                    read_in => sig_read, startOfMachine_out => sig_startOfMachine, reading_out => sig_reading,
                                    type_out => sig_type_out, updateAction_out => sig_updateAction_out, position_out => sig_position_out, size_out => sig_size_out, exp_out => sig_exp_out, man_out => sig_man_out, ready_out => sig_ready_out);


----------------------------------------------------------------------
-- Machine: FASTMem
----------------------------------------------------------------------
------------------------------------
-- Next State Logic (combinatorial)
------------------------------------
FASTMem_NextState: process (mem_counter, FASTByte, sig_read, sig_reading, sig_startOfMachine, FASTMem)
-- machine variables declarations
variable FASTMemory: std_logic_vector(0 to 45111) := X"000B2B31000100010046C001912C56B1236118630F5515E2094C5795815B300AC08201680AFD0379E98080803A535DDF80094C57978080808038303134303630353330B6B3CB80808080808080808080000B2B32000100010047C001912C56B2236118630F5515ED094C5795817B3009C082B1016823DC031FDC8080803A535DEA80094C57978080808038303134313933383638B9B3C080808080808080808080000B2B33000100010046C001912C56B3236118630F551CFE094C5792815B300AC082016D71E803FE8080803A5364FB80094C57978080808038303133383239373830B133B78280808080808080808080000B2B3D000100010048C001912C56BD236118630F6F78F1094C5792815B300AC082016816AB0433FA8080803A6E40ED80094C57978080808038303133383430393336B23338B68280808080808080808080000B2B40000100010048C001912C56C0236118630F7A0FC8094C578E817B3009C082B1016823DC031FDD8080803A7857C380094C57978080808038303133323938383631B532B1B180808080808080808080000B2B47000100010046C001912C56C723611863100D4DEB094C5792815B300AC082016842E71653BD8080803B0C15E680094C57978080808038303134303439333835B1B39980808080808080808080000B2B52000100010047C001912C56D223611863102C24C2094C5792815B300AC082016842F60442B08080803B2A6CBE80094C57978080808038303133393838313035B732B1F180808080808080808080000B2B5D000100010052C001912C56DD23611863103029D5094C579781793C09C080B101681689076DCF0AA380803B2E71D11FA1094C5797094C57973B2E71D28080808038303134323438393939B133B98280808080808080808080000B2B5E000100010051C001912C56DE2361186310302B9F094C579781593C0AC08001680AFD0379EA04A380803B2E739A03F5094C5797094C57973B2E739B8080808038303134323439303030B138B68280808080808080808080000B2B5F000100010052C001912C56DF2361186310302BAA094C579781793C09C080B1016842E71653BE15B580803B2E73A608CD094C5797094C57973B2E73A78080808038303134323439303030B238B6B180808080808080808080000B2B6000010001007DC001912C56E02361186310302CB0094C579783593C0AC080016842E71653BF14D680803B2E74AC0AF9094C5797094C57973B2E74AC8080808038303134323439303030B638B68280808080808080808080218CB48080807AC480808080808680808080808080808080A3C18080808180D0808080808080808080808080000B2B6100010001007EC001912C56E12361186310302E9D094C579783593C0AC080016823DC031FDE019B80803B2E769905BD094C5797094C57973B2E76998080808038303134323439303030B938B68280808080808080808080218CB4FF80808180808080808680808080808080808080A3C18080800111A980D1808080808080808080808080000B2B62000100010051C001912C56E22361186310302F9D094C579781593C0AC080016816AB0433FB0CBC80803B2E77990785094C5797094C57973B2E779A8080808038303134323439303031B238B68280808080808080808080000B2B63000100010052C001912C56E32361186310302FF4094C579781793C09C080B1016816AB0433FC0CD680803B2E77F00785094C5797094C57973B2E77F18080808038303134323439303031B538B68280808080808080808080000B2B64000100010052C001912C56E423611863103033F9094C579781793C09C080B1016842E71653C2158B80803B2E7BF507E9094C5797094C57973B2E7BF58080808038303134323439303031B938B69480808080808080808080000B2B6500010001004FC001912C56E5236118631030348F094C5797815B3C0AC08001682AC86FC2FFA380803B2E7C8B17B9094C5797094C57973B2E7C8C8080808038303134323439303032B0B48B80808080808080808080000B2B6600010001004FC001912C56E623611863103034E2094C5797815B3C0AC08001682AC86FC3FFA280803B2E7CDE17B9094C5797094C57973B2E7CDF8080808038303134323439303032B2B48C80808080808080808080000B2B67000100010050C001912C56E72361186310303591094C579781593C0AC08001682AC86FC4038780803B2E7D8D05BD094C5797094C57973B2E7D8E8080808038303134323439303032B331B08280808080808080808080000B2B68000100010069C001912C56E823611863103035D1094C5797825B3C0AC080016842E71653C3819E80803B2E7DCD02AD094C5797094C57973B2E7DCE8080808038303134323439303032B632B78280808080808080808080238CC180808005BD808080D0808080808080808080808080000B2B69000100010078C001912C56E92361186310303A85094C5792825B300AC082016842F60442B18080803B2F028180094C57978080808038303134303430303034B532B7B080808080808080808080430C0AC080FF00C18080011CA1094C57973B2F02828080808038303134323439303032B932B78980808080808080808080000B2B6A000100010077C001912C56EA2361186310303ADE094C5792825B300AC082016842F60442B38080803B2F02D980094C57978080808038303134303430333235B432B7B180808080808080808080430C0AC080FF00C180802DA9094C57973B2F02DA8080808038303134323439303033B032B78A80808080808080808080000B2B6B000100010051C001912C56EB2361186310303AF6094C579781593C0AC080016823DC031FE1019880803B2F02F200E5094C5797094C57973B2F02F38080808038303134323439303033B132B78380808080808080808080000B2B6C000100010051C001912C56EC2361186310303BD0094C579781593C0AC08001680AFD0379EB049F80803B2F03CC00E5094C5797094C57973B2F03CC8080808038303134323439303033B232B78480808080808080808080000B2B6D000100010077C001912C56ED2361186310303BE8094C5792825B300AC082016842F60442B58080803B2F03E480094C57978080808038303134303430353833B632B7B280808080808080808080430C0AC080FF00C1808021CD094C57973B2F03E58080808038303134323439303033B332B78B80808080808080808080000B2B6E000100010053C001912C56EE2361186310303BF4094C5797817B3C09C080B1016823DC031FE2FF9080803B2F03F001C9094C5797094C57973B2F03F18080808038303134323439303033B43132B98780808080808080808080000B2B6F000100010052C001912C56EF2361186310303FE7094C5797815B3C0AC080016842E71653C5FF028380803B2F07E302AD094C5797094C57973B2F07E48080808038303134323439303033B732B79380808080808080808080000B2B70000100010051C001912C56F02361186310304187094C579781593C0AC08001681689076DD009BC80803B2F098304D9094C5797094C57973B2F09848080808038303134323439303033B837B7AB80808080808080808080000B2B71000100010051C001912C56F12361186310304488094C5797815B3C0AC080016842E71653C6819A80803B2F0C8402AD094C5797094C57973B2F0C848080808038303134323439303034B237B78F80808080808080808080000B2B72000100010050C001912C56F2236118631030479D094C5797815B3C0AC080017423BA5C9AFF01FF80803B2F0F998B094C5797094C57973B2F0F9A8080808038303134323439303034B432B79380808080808080808080000B2B73000100010051C001912C56F323611863103047A4094C5797815B3C0AC08001680AFD0379ECFFB680803B2F0FA008CD094C5797094C57973B2F0FA18080808038303134323439303034B537B78980808080808080808080000B2B74000100010053C001912C56F423611863103048DF094C579781793C09C080B1016842E71653C715E580803B2F10DB21CD094C5797094C57973B2F10DB8080808038303134323439303035B03338B6D380808080808080808080000B2B75000100010051C001912C56F52361186310304A82094C5797815B3C0AC080016842E71653C8819A80803B2F11FE00E5094C5797094C57973B2F11FE8080808038303134323439303035B332B79080808080808080808080000B2B76000100010052C001912C56F62361186310304CBC094C5797817B3C09C080B1017423BA5C9BFF029180803B2F14B8B3094C5797094C57973B2F14B98080808038303134323439303035B83236B28680808080808080808080000B2B77000100010052C001912C56F72361186310304DB2094C579781593C0AC08001680AFD0379ED049680803B2F15AE0CC1094C5797094C57973B2F15AF8080808038303134323439303036B03338B68C80808080808080808080000B2B78000100010053C001912C56F82361186310304DC2094C5797815B3C0AC080016816AB0433FDFF019480803B2F15BE09B1094C5797094C57973B2F15BE8080808038303134323439303036B13338B68780808080808080808080000B2B79000100010051C001912C56F92361186310304EFE094C579781593C0AC080016815F157BC08BF80803B2F16FA04D9094C5797094C57973B2F16FB8080808038303134323439303036B23236B28880808080808080808080000B2B7A000100010053C001912C56FA2361186310304F82094C579781793C09C080B101681689076DD10AB180803B2F16FE00E5094C5797094C57973B2F16FF8080808038303134323439303036B33338B68380808080808080808080000B2B7B000100010052C001912C56FB2361186310304F83094C579781593C0AC08001681689076DD209D380803B2F16FF04D9094C5797094C57973B2F16FF8080808038303134323439303036B43236B2A080808080808080808080000B2B7C000100010052C001912C56FC2361186310304F87094C579781593C0AC080016816AB0433FE0C8680803B2F178303F5094C5797094C57973B2F17848080808038303134323439303036B53236B28580808080808080808080000B2B7D00010001007CC001912C56FD2361186310304F88094C579783793C09C080B1017423BA5C9C14A980803B2F178495094C5797094C57973B2F17858080808038303134323439303036B63338B68280808080808080808080218CB4808080F680808080808680808080808080808080A3C18080808180D1808080808080808080808080000B2B7E000100010053C001912C56FE2361186310304F89094C579781793C09C080B101681689076DD30AF580803B2F178501C9094C5797094C57973B2F17868080808038303134323439303036B73338B6A380808080808080808080000B2B7F000100010053C001912C56FF2361186310304F8F094C5797817B3C09C080B101680AFD0379EEFFB780803B2F178B0FD1094C5797094C57973B2F178C8080808038303134323439303036B83338B68280808080808080808080000B2B80000100010051C001912C578023611863103050C6094C579781593C0AC08001682AC86FC502EE80803B2F18C20EED094C5797094C57973B2F18C28080808038303134323439303037B03236B28880808080808080808080000B2B81000100010052C001912C578123611863103051A5094C579781593C0AC080016843980E3FE1158B80803B2F19A102AD094C5797094C57973B2F19A28080808038303134323439303037B13236B28980808080808080808080000B2B82000100010051C001912C578223611863103052ED094C579781593C0AC08001682AC86FC6038180803B2F1AE914A9094C5797094C57973B2F1AEA8080808038303134323439303037B33236B28380808080808080808080000B2B83000100010051C001912C578323611863103053E0094C579781593C0AC08001680AFD0379EF03A580803B2F1BDC06A1094C5797094C57973B2F1BDD8080808038303134323439303037B432B7DE80808080808080808080000B2B84000100010050C001912C57842361186310305591094C579781593C0AC08001737CED168C058980803B2F1D8D95094C5797094C57973B2F1D8E8080808038303134323439303037B73338B68280808080808080808080000B2B85000100010052C001912C578523611863103055AB094C579781593C0AC080016842E71653C910CA80803B2F1DA701C9094C5797094C57973B2F1DA88080808038303134323439303037B832B701E980808080808080808080000B2B86000100010083C001912C578623611863103062BE094C579783793C09C080B1016842E71653CA14CF80803B2F2ABA024FF9094C5797094C57973B2F2ABB8080808038303134323439303038B13236B28380808080808080808080218CB48080807D3DAC80808080808680808080808080808080A3C180808002369580D1808080808080808080808080000B2B87000100010053C001912C578723611863103075FA094C5797817B3C09C080B1016842F60442B7FF00C780803B2F3DF607E9094C5797094C57973B2F3DF78080808038303134323439303038B739B8A680808080808080808080000B2B88000100010051C001912C57882361186310307689094C579781593C0AC080016842E71653CD14B480803B2F3E8500E5094C5797094C57973B2F3E868080808038303134323439303038B839B88480808080808080808080000B2B89000100010052C001912C578923611863103076F6094C579781793C09C080B101680AFD0379F004B580803B2F3EF203F5094C5797094C57973B2F3EF38080808038303134323439303038B939B88580808080808080808080000B2B8A000100010053C001912C578A2361186310307788094C579781793C09C080B101680AFD0379F104C380803B2F3F840058A5094C5797094C57973B2F3F858080808038303134323439303039B039B88980808080808080808080000B2B8B000100010051C001912C578B2361186310307796094C579781593C0AC080016842F60442B8059280803B2F3F9203F5094C5797094C57973B2F3F938080808038303134323439303039B139B88280808080808080808080000B2B8C000100010051C001912C578C23611863103077F3094C5797817B3C09C080B1016D71E803FFFF00F780803B2F3FEF9F094C5797094C57973B2F3FF08080808038303134323439303039B239B88280808080808080808080000B2B8D000100010050C001912C578D23611863103078B2094C579781793C09C080B101737CED168D05D180803B2F40AE8E094C5797094C57973B2F40AF8080808038303134323439303039B339B88480808080808080808080000B2B8E000100010050C001912C578E23611863103078C1094C5797817B3C09C080B1017040900699818280803B2F40BD90094C5797094C57973B2F40BE8080808038303134323439303039B439B88680808080808080808080000B2B8F000100010054C001912C578F236118631030798E094C5797817B3C09C080B1016842E71653CEFF02BB80803B2F418A17B9094C5797094C57973B2F418A8080808038303134323439303039B537B702D480808080808080808080000B2B9000010001004FC001912C57902361186310307ACB094C579781593C0AC080016D738D25B00A8580803B2F42C798094C5797094C57973B2F42C88080808038303134323439303039B639B88380808080808080808080";

begin
	NextState_FASTMem <= FASTMem;
	-- Set default values for outputs and signals
	sig_read <= '1';
    next_sig_msg_in <= sig_msg_in;
	next_mem_counter <= mem_counter;
	case FASTMem is
		when Start =>
			IF (sig_startOfMachine = '1' AND sig_reading = '0') THEN
				sig_read <= '1';
			ELSIF (sig_startOfMachine = '0' AND sig_reading = '1') THEN
				sig_read <= '1';
			ELSIF (sig_startOfMAchine = '0' AND sig_reading = '0') THEN
				sig_read <= '0';
			END IF;
			if sig_read = '1' then
				NextState_FASTMem <= writeByte;
			end if;
		when writeByte =>
			IF (sig_reading = '1') THEN
				next_sig_msg_in <= FASTMemory(mem_counter to (mem_counter + 7));
				next_mem_counter <= mem_counter + 8;
			END IF;
			if sig_startOfMachine = '1' then
				NextState_FASTMem <= Start;
			else
				NextState_FASTMem <= writeByte;
			end if;
--vhdl_cover_off
		when others =>
			null;
--vhdl_cover_on
	end case;
end process;

------------------------------------
-- Current State Logic (sequential)
------------------------------------
FASTMem_CurrentState: process (sig_clk)
begin
	if rising_edge(sig_clk) then
		if sig_reset = '1' then
			FASTMem <= Start;
		else
			if sig_enable = '1' then
				FASTMem <= NextState_FASTMem;
			end if;
		end if;
	end if;
end process;

------------------------------------
-- Registered Outputs Logic
------------------------------------
FASTMem_RegOutput: process (sig_clk)
begin
	if rising_edge(sig_clk) then
		if sig_reset = '1' then
			-- FASTByte <= 		-- Initialization in the reset state or default value required!
			-- mem_counter <= 		-- Initialization in the reset state or default value required!
		else
			if sig_enable = '1' then
				sig_msg_in <= next_sig_msg_in;
				mem_counter <= next_mem_counter;
			end if;
		end if;
	end if;
end process;

bookHandler: process (sig_clk)
begin
    if rising_edge(sig_clk) then
		if sig_reset = '1' then

            counter <= 0;

            bidOrderDepthBook_size <= (OTHERS => X"0000000000000000");
            bidOrderDepthBook_px_exp <= (OTHERS => X"00000000");
            bidOrderDepthBook_px_man <= (OTHERS => X"FFFFFFFFFFFFFFFF");

            offerOrderDepthBook_size <= (OTHERS => X"0000000000000000");
            offerOrderDepthBook_px_exp <= (OTHERS => X"00000000");
            offerOrderDepthBook_px_man  <= (OTHERS => X"FFFFFFFFFFFFFFFF");
		else
			if sig_enable = '1' then

                counter <= counter + 1;

				--
                IF (sig_ready_out = '1') THEN
                    IF (sig_type_out = '0') THEN			-- bid
                            
                        for i in 9 downto 1 loop		                                        -- position shift (testar depois pq coloquei 1 agora, tava 0)
                            bidOrderDepthBook_size(i) <= bidOrderDepthBook_size(i - 1);
                            bidOrderDepthBook_px_exp(i) <= bidOrderDepthBook_px_exp(i - 1);
                            bidOrderDepthBook_px_man(i) <= bidOrderDepthBook_px_man(i - 1);
                            if i = to_integer(unsigned(sig_position_out)) then
                                    exit;
                            end if;
                        end loop;

                        bidOrderDepthBook_size(to_integer(signed(sig_position_out - 1))) <= sig_size_out;
                        bidOrderDepthBook_px_exp(to_integer(signed(sig_position_out - 1))) <= sig_exp_out;
                        bidOrderDepthBook_px_man(to_integer(signed(sig_position_out - 1))) <= sig_man_out;

                    ELSIF (sig_type_out = '1') THEN		-- offer
                    
                        for i in 9 downto 1 loop                                        		-- position shift
                            offerOrderDepthBook_size(i) <= offerOrderDepthBook_size(i - 1);
                            offerOrderDepthBook_px_exp(i) <= offerOrderDepthBook_px_exp(i - 1);
                            offerOrderDepthBook_px_man(i) <= offerOrderDepthBook_px_man(i - 1);
                            if i = to_integer(unsigned(sig_position_out)) then
                                    exit;
                            end if;
                        end loop;

                        offerOrderDepthBook_size(to_integer(signed(sig_position_out - 1))) <= sig_size_out;
                        offerOrderDepthBook_px_exp(to_integer(signed(sig_position_out - 1))) <= sig_exp_out;
                        offerOrderDepthBook_px_man(to_integer(signed(sig_position_out - 1))) <= sig_man_out;
                    END IF;
                END IF;
                --
			end if;
		end if;
	end if;
end process;



END ARCHITECTURE;
